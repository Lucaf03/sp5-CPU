library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package sp_pkg is

  type INSTR_NAME is (
    ADD, SUB, SLLR, SLT, SLTU, XORR, SRLR, SRAR, ORR, ANDR,
    ADDI, SLTI, SLTIU, XORI, ORI, ANDI, SLLI, SRLI, SRAI,
    LB, LH, LW, LBU, LHU,
    SB, SH, SW,
    BEQ, BNE, BLT, BGE, BLTU, BGEU,
    LUI, AUIPC,
    JAL, JALR,
    NOP,
    MUL, MULH, MULHSU, MULHU, DIV, DIVU, REMM, REMU,
    CSRRW, CSRRS, CSRRC, CSRRWI, CSRRSI, CSRRCI
  );

  constant mvendorid_addr : std_logic_vector(11 downto 0)  := x"F11";
  constant marchid_addr : std_logic_vector(11 downto 0)   := x"F12";
  constant mimpid_addr : std_logic_vector(11 downto 0)    := x"F13";
  constant mhartid_addr : std_logic_vector(11 downto 0)   := x"F14";
  constant mstatus_addr : std_logic_vector(11 downto 0)   := x"300";
  constant misa_addr : std_logic_vector(11 downto 0)      := x"301";

end package sp_pkg;
